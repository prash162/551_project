module sll_slh(offset,SreadA,sll_slh_out);
  input [15:0] offset;
  input [15:0] SreadA;
  output [15:0]sll_slh_out;
endmodule
