
module decoder(Instr, VADD,VDOT,SMUL,SST,VLD,VST,SLL,SLH,J,NOP);
input [3:0] Instr; 
output VADD,VDOT,SMUL,SST,VLD,VST,SLL,SLH,J,NOP;

reg VADD,VDOT,SMUL,SST,VLD,VST,SLL,SLH,J,NOP;

always@(Instr)
begin
	case(Instr)	
		4'b0000:
			{VADD,VDOT,SMUL,SST,VLD,VST,SLL,SLH,J,NOP} = 10'b1000000000;
		4'b0001:
			{VADD,VDOT,SMUL,SST,VLD,VST,SLL,SLH,J,NOP} = 10'b0100000000;
		4'b0010:
			{VADD,VDOT,SMUL,SST,VLD,VST,SLL,SLH,J,NOP} = 10'b0010000000;
		4'b0011:
			{VADD,VDOT,SMUL,SST,VLD,VST,SLL,SLH,J,NOP} = 10'b0001000000;
		4'b0100:
			{VADD,VDOT,SMUL,SST,VLD,VST,SLL,SLH,J,NOP} = 10'b0000100000;
		4'b0101:
			{VADD,VDOT,SMUL,SST,VLD,VST,SLL,SLH,J,NOP} = 10'b0000010000;
		4'b0110:
			{VADD,VDOT,SMUL,SST,VLD,VST,SLL,SLH,J,NOP} = 10'b0000001000;
		4'b0111:
			{VADD,VDOT,SMUL,SST,VLD,VST,SLL,SLH,J,NOP} = 10'b0000000100;
		4'b1000:
			{VADD,VDOT,SMUL,SST,VLD,VST,SLL,SLH,J,NOP} = 10'b0000000010;
		4'b1111:
			{VADD,VDOT,SMUL,SST,VLD,VST,SLL,SLH,J,NOP} = 10'b0000000001;
		default:
			{VADD,VDOT,SMUL,SST,VLD,VST,SLL,SLH,J,NOP} = 10'b0000000000;

	

	endcase
end
endmodule
