module sll_slh(offset,SreadA,sll_slh_out);
endmodule
